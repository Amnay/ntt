
program automatic test;

    Environment env;
    initial begin
        env.new();
        env.build();
        env.run();
    end

endprogram
